import uvm_pkg::*;
`include "uvm_macros.svh"

class risc_env extends uvm_env;
    `uvm_component_utils(risc_env)

    risc_agent    agent;
    risc_coverage  coverage;
    risc_scoreboard scoreboard;

    function new(string name = "risc_env", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        agent     = risc_agent::type_id::create("agent", this);
        coverage  = risc_coverage::type_id::create("coverage", this);
        scoreboard = risc_scoreboard::type_id::create("scoreboard", this);
    endfunction

    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        agent.monitor.instr_inport.connect(coverage.analysis_export);
        agent.monitor.memory_inport.connect(scoreboard.memory_export);
    endfunction
endclass
